module spi_master(
// SPI master with proper 8-bit transfer (Mode 0, SCLK idle low)
    input clk,
    input rst,
    input [7:0] data_in,
    input start,
    output reg sclk,
    output reg mosi,
    output reg cs,
    output reg done
);
    reg [3:0] bit_cnt;
    reg [7:0] shift_reg;
    reg [1:0] state;
    localparam IDLE=0, LOAD=1, TRANSFER=2, FINISH=3;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            sclk <= 0; // Mode 0: idle low
            mosi <= 0;
            cs   <= 1;
            done <= 0;
            bit_cnt <= 0;
            shift_reg <= 0;
        end else begin
            case(state)
                IDLE: begin
                    sclk <= 0;
                    cs <= 1;
                    done <= 0;
                    if (start) begin
                        cs <= 0;
                        shift_reg <= data_in;
                        bit_cnt <= 4'd7;
                        state <= LOAD;
                    end
                end
                LOAD: begin
                    mosi <= shift_reg[7];
                    state <= TRANSFER;
                end
                TRANSFER: begin
                    sclk <= 1;
                    state <= FINISH;
                end
                FINISH: begin
                    sclk <= 0;
                    shift_reg <= {shift_reg[6:0],1'b0};
                    if (bit_cnt == 0) begin
                        cs <= 1;
                        done <= 1;
                        state <= IDLE;
                    end else begin
                        bit_cnt <= bit_cnt - 1;
                        state <= LOAD;
                    end
                end
            endcase
        end
    end
endmodule
